interface adder_if();
    logic clk; 
    logic [7:0] a;
    logic [7:0] b;
    logic [8:0] y;
endinterface

`include "uvm_macros.svh"
import uvm_pkg::*; // 전체 라이브러리 전부 끌어오기

class adder_seq_item extends uvm_sequence_item;
    rand bit [7:0] a;
    rand bit [7:0] b;
    bit [8:0] y;
    function new(string name = "ADDER_ITEM");
        super.new(name);
    endfunction

    `uvm_object_utils_begin(adder_seq_item)
        `uvm_field_int(a,UVM_DEFAULT) 
        `uvm_field_int(b,UVM_DEFAULT)
        `uvm_field_int(y,UVM_DEFAULT)
    `uvm_object_utils_end
endclass

class adder_sequence extends uvm_sequence #(adder_seq_item);
    `uvm_object_utils(adder_sequence)
    function new(string name = "SEQ"); //component 상속 ㄴㄴ
        super.new(name);
    endfunction

    adder_seq_item adder_item;

    virtual task body(); //phase 단위 ㄴㄴ
        adder_item = adder_seq_item::type_id::create("ADDER_ITEM");
        for(int i=0; i<10; i++) begin
            start_item(adder_item);
            adder_item.randomize();
            `uvm_info("SEQ",$sformatf("adder item to driver a:%0d,b:%0d",adder_item.a,adder_item.b),UVM_NONE)
            adder_item.print(uvm_default_line_printer);

            finish_item(adder_item);


        end
    endtask //s
endclass
class adder_driver extends uvm_driver #(adder_seq_item);
    `uvm_component_utils(adder_driver)
    function new(string name = "DRV", uvm_component parent);
       super.new(name,parent);
    endfunction //new()

    adder_seq_item adder_item;
    virtual adder_if a_if;

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        adder_item = adder_seq_item::type_id::create("ADDER_ITEM");

        if(!uvm_config_db#(virtual adder_if)::get(this,"","a_if",a_if))
            `uvm_fatal("DRV","adder_if not found via uvm_config_db")
    endfunction

    virtual task run_phase(uvm_phase phase);
        
        forever begin
            seq_item_port.get_next_item(adder_item);
            @(posedge a_if.clk);
            a_if.a = adder_item.a;
            a_if.b = adder_item.b;
            

            `uvm_info("DRV",$sformatf("DRIVE DUT a:%0d,b:%0d",adder_item.a,adder_item.b),UVM_LOW)
            adder_item.print(uvm_default_line_printer);

            seq_item_port.item_done();
            // #10;
        end

    endtask
endclass //adder_driver 

class adder_monitor extends uvm_monitor;    
    `uvm_component_utils(adder_monitor)
    uvm_analysis_port #(adder_seq_item) send; 
    function new(string name = "MON", uvm_component parent);
        super.new(name, parent);
        send = new("WRITE", this);
    endfunction //new()

    adder_seq_item adder_item;
    virtual adder_if a_if;

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase); // item 생성 
        adder_item = adder_seq_item::type_id::create("ADDER_ITEM"); //연결
        if(!uvm_config_db#(virtual adder_if)::get(this,"","a_if",a_if)) 
            `uvm_fatal("MON","adder_if not found in uvm_config_db")
    endfunction

    virtual task run_phase(uvm_phase phase);
   
       forever begi 알아서 analysis_port에 연결 // ㅁㅁㅁㅁㅎscoreㅂ보볻보보보드등드드드으의의의의 recive ㅇ여연연연연ㄱ겨결결결결n
            // #10;
            @(posedge a_if.clk);
            #1;
            adder_item.a = a_if.a;
            adder_item.b = a_if.b;
            adder_item.y = a_if.y;

           `uvm_info("MON",$sformatf("sampled a: %0d,b:%0d,y:%0d",adder_item.a,adder_item.b,adder_item.y),UVM_LOW)
           adder_item.print(uvm_default_line_printer);

           send.write(adder_item); //send to scb  알아서 analysis_port에 연결 
       end 
    endtask //



endclass //adder_monitor
class adder_scoreboard extends uvm_scoreboard;
    `uvm_component_utils(adder_scoreboard) // factory 등록

    uvm_analysis_imp #(adder_seq_item,adder_scoreboard) recv; // uvm 제공 class recv:핸들러
    adder_seq_item adder_item; // tranaction 받기

    function new(string name = "SCO", uvm_component parent);
        super.new(name,parent);
        recv = new("READ", this);
    endfunction //new()

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        adder_item = adder_seq_item::type_id::create("ADDER_ITEM");
    endfunction

    virtual function void write(adder_seq_item item); //transaction 값 저장 
        adder_item = item;
        `uvm_info("SCO",$sformatf("Receive a:%0d, b:%0d, y:%0d",item.a,item.b,item.y),UVM_LOW)
        adder_item.print(uvm_default_line_printer);

        if(adder_item.y == adder_item.a + adder_item.b)
            `uvm_info("SCO","*** TEST PASSED ***",UVM_NONE)
        else
            `uvm_error("SCO","*** TEST FAILD ***")
    endfunction

endclass //adder_scoreboar

class adder_agent extends uvm_agent;
    `uvm_component_utils(adder_agent) // factory 등록
    function new(string name = "AGENT", uvm_component parent);
        super.new(name,parent);    
    endfunction

    adder_monitor adder_mon;
    adder_driver adder_drv;
    uvm_sequencer #(adder_seq_item) adder_sqr; //sequncer는 내장된 클래스 사용

    virtual function void build_phase(uvm_phase phase);
       super.build_phase(phase);
       adder_mon = adder_monitor::type_id::create("MON",this);
       adder_drv = adder_driver::type_id::create("DRV",this);
       adder_sqr = uvm_sequencer#(adder_seq_item)::type_id::create("SQR",this);        
    endfunction 

    virtual function void connect_phase(uvm_phase phase);
       super.connect_phase(phase);
       adder_drv.seq_item_port.connect(adder_sqr.seq_item_export); // port와 export 연결 
    endfunction
endclass

class adder_envirnment extends uvm_env;
    `uvm_component_utils(adder_envirnment) //factory에 등록

    function new(string name = "ENV", uvm_component parent);
        super.new(name,parent); 
    endfunction

    adder_scoreboard adder_sco; 알아서 analysis_port에 연결 // ㅁㅁㅁㅁㅎscoreㅂ보볻보보보드등드드드으의의의의 recive ㅇ여연연연연ㄱ겨결결결결
    adder_agent adder_agt;

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        adder_sco = adder_scoreboard::type_id::create("SCO",this);
        adder_agt = adder_agent::type_id::create("AGT",this);
    endfunction

    virtual function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);// 
        adder_agt.adder_mon.send.connect(adder_sco.recv);  // TLM Port와 연결 // score보드의 recive 연결
        
    endfunction
endclass


class test extends uvm_test; //uvm library에 있는거 그대로 상속 // 접근한다고 생각 
    `uvm_component_utils(test) //factory에 등록 매크로 
    function new(string name = "TEST", uvm_component parent); 
        super.new(name,parent); //super:부모 클래스 

    endfunction //new()
    adder_sequence adder_seq;
    adder_envirnment adder_env; //handler

    virtual function void build_phase(uvm_phase phase); // uvm에서 제공해주는 클래스이름 component에 있음
        super.build_phase(phase);
        adder_seq = adder_sequence::type_id::create("SEQ",this); //factory excute
        adder_env = adder_envirnment::type_id::create("ENV",this); // sysverilog의 new랑 비슷 
    endfunction 
    //sequencer : generator 느낌임 sequence: transaction 느낌
    virtual task run_phase(uvm_phase phase); // 함수 구현 : override 하기  
        phase.raise_objection(phase); //drop전까지 simulation이 끝나지 않는다. 
        adder_seq.start(adder_env.adder_agt.adder_sqr); //sequence랑 sequencer랑 다름
        phase.drop_objection(phase); //objection 해제. run_phase 
    endtask 

endclass //test ext

module tb_adder();
    test adder_test;
    adder_if a_if();

    adder dut(
        .a(a_if.a),
        .b(a_if.b),
        .y(a_if.y)
    );
always #5 a_if.clk = ~a_if.clk;
initial begin
    a_if.clk = 0;
    adder_test = new("TEST",null);
    uvm_config_db #(virtual adder_if)::set(null, "*","adder_if",a_if); // interface에 대한 정보 저장 db에
   
    run_test();

end

endmodule
